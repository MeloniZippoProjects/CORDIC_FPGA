library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library cordic;

use cordic.util.all;

entity atan_lut_15x32 is
	port (
		iteration	: in	std_ulogic_vector (f_log2(15)-1 downto 0);
		atan		: out	std_ulogic_vector (31 downto 0)
	);
end atan_lut_15x32;

architecture rtl of atan_lut_15x32 is

	signal addr_int 	: integer range 0 to 14;
	type lut_t is array (0 to 14) of std_ulogic_vector (31 downto 0);
	constant lut : lut_t :=
	("00011101101011000110011100000101", "00001111101011011011101011111100", "00000111111101010110111010100110", "00000011111111101010101101110110", "00000001111111111101010101011011", "00000000111111111111101010101010", "00000000011111111111111101010101", "00000000001111111111111111101010", "00000000000111111111111111111101", "00000000000011111111111111111111", "00000000000001111111111111111111", "00000000000000111111111111111111", "00000000000000011111111111111111", "00000000000000001111111111111111", 
	"00000000000000000111111111111111"
	);

	
begin
	addr_int <= TO_INTEGER(unsigned(iteration));
	atan <= lut(addr_int);
end rtl;